`timescale 1ns/10ps
module decoder5_32(in, out, en);

input [4:0] in;
input en;
output [31:0] out;

wire [3:0] dec24_out;

decoder2_4 dec24 (in[4:3], dec24_out, en);

decoder3_8 dec38_0 (in[2:0], out[7:0], dec24_out[0]);
decoder3_8 dec38_1 (in[2:0], out[15:8], dec24_out[1]);
decoder3_8 dec38_2 (in[2:0], out[23:16], dec24_out[2]);
decoder3_8 dec38_3 (in[2:0], out[31:24], dec24_out[3]);

endmodule


module decoder_5to32_test;
reg [4:0] in;
reg en;
wire [31:0] out;

decoder5_32 test (.in, .out, .en);

initial begin
	en = 1;
	in = 5'b00000; #500;
	in = 5'b00001; #500;
	in = 5'b00010; #500;
	in = 5'b00011; #500;
	in = 5'b00100; #500;
	in = 5'b00101; #500;
	in = 5'b00110; #500;
	in = 5'b00111; #500;
	in = 5'b01000; #500;
	in = 5'b01001; #500;
	in = 5'b01011; #500;
	in = 5'b01100; #500;
	in = 5'b01101; #500;
	in = 5'b01110; #500;
	in = 5'b01111; #500;
	in = 5'b10000; #500;
	in = 5'b10001; #500;
	in = 5'b10010; #500;
	in = 5'b10011; #500;
	in = 5'b10100; #500;
	in = 5'b10101; #500;
	in = 5'b10110; #500;
	in = 5'b10111; #500;
	in = 5'b11000; #500;
	in = 5'b11001; #500;
	in = 5'b11010; #500;
	in = 5'b11011; #500;
	in = 5'b11100; #500;
	in = 5'b11101; #500;
	in = 5'b11110; #500;
	in = 5'b11111; #500;
	
	in = 5'b00000; #500;
	in = 5'b00001; #500;
	in = 5'b00010; #500;
	in = 5'b00011; #500;
	in = 5'b00100; #500;
	in = 5'b00101; #500;
	in = 5'b00110; #500;
	in = 5'b00111; #500;
	in = 5'b01000; #500;
	in = 5'b01001; #500;
	in = 5'b01011; #500;
	in = 5'b01100; #500;
	in = 5'b01101; #500;
	in = 5'b01110; #500;
	in = 5'b01111; #500;
	in = 5'b10000; #500;
	in = 5'b10001; #500;
	in = 5'b10010; #500;
	in = 5'b10011; #500;
	in = 5'b10100; #500;
	in = 5'b10101; #500;
	in = 5'b10110; #500;
	in = 5'b10111; #500;
	in = 5'b11000; #500;
	in = 5'b11001; #500;
	in = 5'b11010; #500;
	in = 5'b11011; #500;
	in = 5'b11100; #500;
	in = 5'b11101; #500;
	in = 5'b11110; #500;
	in = 5'b11111; #500;
	
	en = 0;
	in = 5'b00000; #500;
	in = 5'b00001; #500;
	in = 5'b00010; #500;
	in = 5'b00011; #500;
	in = 5'b00100; #500;
	in = 5'b00101; #500;
	in = 5'b00110; #500;
	in = 5'b00111; #500;
	in = 5'b01000; #500;
	in = 5'b01001; #500;
	in = 5'b01011; #500;
	in = 5'b01100; #500;
	in = 5'b01101; #500;
	in = 5'b01110; #500;
	in = 5'b01111; #500;
	in = 5'b10000; #500;
	in = 5'b10001; #500;
	in = 5'b10010; #500;
	in = 5'b10011; #500;
	in = 5'b10100; #500;
	in = 5'b10101; #500;
	in = 5'b10110; #500;
	in = 5'b10111; #500;
	in = 5'b11000; #500;
	in = 5'b11001; #500;
	in = 5'b11010; #500;
	in = 5'b11011; #500;
	in = 5'b11100; #500;
	in = 5'b11101; #500;
	in = 5'b11110; #500;
	in = 5'b11111; #500;

 end

endmodule